// The cumulative top level module for the ECE 271 final project.
// device_switch: A switch which toggles between the nes and ps2
//                controllers. 0 is nes, 1 is ps2.
// reset: Brings the device to its initalization state. This should
//        start on and then be turned off.
// vcc: Used for some protocols.
// gnd: Used for some protocols.
// sys_clk: a 50MHz clock.
// hex1: A number formatted for a hexidecimal 7segment display. It is
//       the least significant digit. It is determind by the current
//       active driver's input.
// hex2: Ibid, but for the most significant digit.
// ps2_data: Pin as per ps2 device protocl.
// CLK_K: Clock generated by the ps2 device.
module g21_final(input logic device_switch, input logic reset, output logic vcc, output logic gnd, //Generic system controls
	input logic sys_clk//VGA driver
	output logic[6:0] hex1, output logic[6:0] hex2,//7seg outputs
	input logic ps2_data, inout logic CLK_K //PS2 pins
	); //NES inputs
	assign vcc 1;
	assign gnd 0;
	
	logic [7:0] ps2_key;
	logic [3:0] nes_key; /*I don't actually know how long your NES key is, but
	it doesn't matter. It can be truncated or modulus'd into the mux, and if
	it is any shorter, it does NOT need to be inflated to 8 bits. The hash 
	function can take smaller values.*/
	logic [7:0] live_key; /*This is the key which is driving the 7seg and VGA.
	At any given point, it will be ps2_key or nes_key*/
	
	
	assign nes_k = 4b'1111; //TODO: REPLACE THIS WITH THE NES DRIVER.
	listener_ps2 ps2_driver(.block(reset), .data(ps2_data), .CLK_K(CLK_K), .key(key));
	
	/*Simple mux: */
	always_comb begin
		if(device_switch) begin //1: PS2
			live_key = ps2_key;
		end else begin
			live_key = nes_key;
		end
	end
	
	/* Output 1: 7seg */
	//None of our devices will give us a big hexidecimal number. Only 2 7segs are needed.
	logic[2:0][3:0] hexidecimal;
	hex_notation splitter #(INPUT_SIZE = 8) (.number(live_key),.hex(hexidecimal));
	sevenseg printer1 (.data(hexidecimal[0]),.segments(hex1));
	sevenseg printer2 (.data(hexidecimal[1]),.segments(hex2));
	
	/* Output 2: RGB */
	logic [31:0] hash;
	chash ec(live_key, hash);
	monitor vga(.reset(reset), .sys_clk(sys_clk), .c_switches(hash%(2**5)),
	.hsync(hsync), .vsync(vsync), .red(red), .green(green), .blue(blue));
endmodule

/* From lab 6:
module monitor
(input logic reset, input logic sys_clk, input logic[5:0] c_switches, 
output logic hsync, output logic vsync, 
output logic [3:0] red, output logic [3:0] green, output logic[3:0] blue);
*/